netcdf simple_nc4 {
dimensions:
	x = 6 ;
	y = 12 ;

group: grp1 {
  variables:
  	uint64 data(x, y) ;
  data:

   data =
  0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11,
  12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23,
  24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35,
  36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47,
  48, 49, 50, 51, 52, 53, 54, 55, 56, 57, 58, 59,
  60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71 ;
  } // group grp1

group: grp2 {
  types:
    compound sample_compound_type {
      int i1 ;
      int i2 ;
    }; // sample_compound_type
  variables:
  	sample_compound_type data(x, y) ;
  data:

   data =
  {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42}, 
      {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42},
  {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42}, 
      {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42},
  {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42}, 
      {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42},
  {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42}, 
      {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42},
  {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42}, 
      {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42},
  {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42}, 
      {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42}, {42, -42} ;
  } // group grp2
}
